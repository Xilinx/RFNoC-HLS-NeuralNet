`timescale 1ns/1ps
`define NS_PER_TICK 1
`define NUM_TEST_CASES 4

`include "sim_exec_report.vh"
`include "sim_clks_rsts.vh"
`include "sim_rfnoc_lib.svh"

module noc_block_ex1layer_tb();
  `TEST_BENCH_INIT("noc_block_ex1layer",`NUM_TEST_CASES,`NS_PER_TICK);
  localparam BUS_CLK_PERIOD = $ceil(1e9/166.67e6);
  localparam CE_CLK_PERIOD  = $ceil(1e9/200e6);
  localparam NUM_CE         = 1;  // Number of Computation Engines / User RFNoC blocks to simulate
  localparam NUM_STREAMS    = 1;  // Number of test bench streams
  `RFNOC_SIM_INIT(NUM_CE, NUM_STREAMS, BUS_CLK_PERIOD, CE_CLK_PERIOD);
  `RFNOC_ADD_BLOCK(noc_block_ex1layer, 0);

  localparam SPP = 784; // Samples per packet

  /********************************************************
  ** Verification
  ********************************************************/
  initial begin : tb_main
    string s;
    logic [31:0] random_word;
    logic [63:0] readback;
    integer data_file; // file handler
    integer scan_file; // file handler

    /********************************************************
    ** Test 1 -- Reset
    ********************************************************/
    `TEST_CASE_START("Wait for Reset");
    while (bus_rst) @(posedge bus_clk);
    while (ce_rst) @(posedge ce_clk);
    `TEST_CASE_DONE(~bus_rst & ~ce_rst);

    /********************************************************
    ** Test 2 -- Check for correct NoC IDs
    ********************************************************/
    `TEST_CASE_START("Check NoC ID");
    // Read NOC IDs
    tb_streamer.read_reg(sid_noc_block_ex1layer, RB_NOC_ID, readback);
    $display("Read EX1LAYER NOC ID: %16x", readback);
    `ASSERT_ERROR(readback == noc_block_ex1layer.NOC_ID, "Incorrect NOC ID");
    `TEST_CASE_DONE(1);

    /********************************************************
    ** Test 3 -- Connect RFNoC blocks
    ********************************************************/
    `TEST_CASE_START("Connect RFNoC blocks");
    `RFNOC_CONNECT(noc_block_tb,noc_block_ex1layer,S16,SPP);
    `RFNOC_CONNECT(noc_block_ex1layer,noc_block_tb,S16,SPP);
    `TEST_CASE_DONE(1);

    /********************************************************
    ** Test 4 -- Write / readback user registers
    ********************************************************/
    `TEST_CASE_START("Write / readback user registers");
    tb_streamer.write_user_reg(sid_noc_block_ex1layer, noc_block_ex1layer.SR_SIZE_INPUT, SPP*4);
    tb_streamer.read_user_reg(sid_noc_block_ex1layer, noc_block_ex1layer.RB_SIZE_INPUT, readback);
    $sformat(s, "User register 0 incorrect readback! Expected: %0d, Actual %0d", readback[31:0], SPP*4);
    `ASSERT_ERROR(readback[31:0] == SPP*4, s);
    random_word = $random();
    tb_streamer.write_user_reg(sid_noc_block_ex1layer, noc_block_ex1layer.SR_SIZE_OUTPUT, 10*4);
    tb_streamer.read_user_reg(sid_noc_block_ex1layer, noc_block_ex1layer.RB_SIZE_OUTPUT, readback);
    $sformat(s, "User register 1 incorrect readback! Expected: %0d, Actual %0d", readback[31:0], 10*4);
    `ASSERT_ERROR(readback[31:0] == 10*4, s);
    `TEST_CASE_DONE(1);

    /********************************************************
    ** Test 5 -- Test sequence
    ********************************************************/
    // ex1layer's user code is a loopback, so we should receive
    // back exactly what we send
    // `TEST_CASE_START("Test sequence");
    // fork
    //   begin
    //     cvita_payload_t send_payload;
    //     for (int i = 0; i < SPP/2; i++) begin
    //       send_payload.push_back(64'(i));
    //     end
    //     tb_streamer.send(send_payload);
    //   end
    //   begin
    //     cvita_payload_t recv_payload;
    //     cvita_metadata_t md;
    //     logic [63:0] expected_value;
    //     tb_streamer.recv(recv_payload,md);
    //     for (int i = 0; i < SPP/2; i++) begin
    //       expected_value = i;
    //       $sformat(s, "Incorrect value received! Expected: %0d, Received: %0d", expected_value, recv_payload[i]);
    //       `ASSERT_ERROR(recv_payload[i] == expected_value, s);
    //     end
    //   end
    // join
    // `TEST_CASE_DONE(1);


    fork
      begin
        real data_float;
        integer data_int;
        logic [15:0] data_logic;
        data_file = $fopen("mnist_validation_data_784x1.dat", "r");
        `ASSERT_FATAL(data_file != 0, "Data file could not be opened");
        if (data_file == 0) begin
          $display("data_file handle was NULL");
          $finish;
        end
        $display("Send data from text file");
        while (!$feof(data_file)) begin
          scan_file = $fscanf(data_file, "%f", data_float);
          data_int = data_float * (2**10);
          data_logic = data_int;
          if (!$feof(data_file))
            tb_streamer.push_word({data_logic}, 0 );
          else
            tb_streamer.push_word({data_logic}, 1 );
          $sformat(s, "Pushing word: %f, %d", data_float, data_int);
          //$display(s);
        end
        $fclose(data_file);
      end
      begin
        logic last;
        logic [15:0] res_logic;
        shortint res_int;
        real res_float;
        // logic [15:0] idx_ref, mag_ref;
        // integer idx_samp_int, mag_samp_int, idx_ref_int, mag_ref_int;
        // $display("Receive FIR filter output");
        // data_file_ref = $fopen("../../../../data_ref_gmsk.txt", "r");
        // `ASSERT_FATAL(data_file_ref != 0, "Output data file could not be opened");
        // data_file_out = $fopen("../../../../data_out_gmsk.txt", "w");
        // `ASSERT_FATAL(data_file_out != 0, "Output data file could not be opened");
        // last = 0;
        for (int ii = 0; ii < 10; ii++) begin
          tb_streamer.pull_word({res_logic}, last);
          res_int = res_logic;
          res_float =  res_int / 2.0**8;
          $sformat(s, "Received Value: %f", res_float);
          $display(s);
          // scan_file = $fscanf(data_file_ref, "%d %d\n", idx_ref, mag_ref);
          // idx_samp_int = idx_samp; mag_samp_int = mag_samp;
          // idx_ref_int = idx_ref;   mag_ref_int = mag_ref;
          // // Check I / Q values, should be equivalent to reference
          // $sformat(s, "Incorrect output value received! Expected: %0d, %0d Received: %0d, %0d", idx_ref_int, mag_ref_int, idx_samp_int, mag_samp_int);
          // `ASSERT_ERROR((mag_samp_int - mag_ref_int) < 50 && (mag_ref_int-mag_samp_int) > -50, s);
          // $fwrite(data_file_out,"%d %d\n", idx_samp, mag_samp);
        end
        // $fclose(data_file_ref);
        // $fclose(data_file_out);
      end
    join
    `TEST_CASE_DONE(1);


    `TEST_BENCH_DONE;

  end
endmodule
